library IEEE;
	use IEEE.STD_LOGIC_1164.all;
	use IEEE.NUMERIC_STD.ALL;

package FIR_Filter_2_package is

constant input_width : positive := 24;
constant output_width : positive := 24;
constant taps : positive := 128;
constant coefficient_width :positive:= 16;

type coefficient_array is array(0 to (taps/2)-1) of signed(coefficient_width-1 downto 0);
constant coefficient : coefficient_array := (
"1000000000000000","1000000000000000","1000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","1000000000000000",
"1000000000000010","1000000000000010","0000000000000000","0000000000000111","0000000000001110","0000000000001010","1000000000010000","1000000000110111",
"1000000001000100","1000000000001000","0000000010000100","0000000100000010","0000000011000101","1000000010011110","1000001010001111","1000001101001001",
"1000000011110010","0000010001001010","0000100001110001","0000011101100111","1000001011010010","1000110000111110","1000110110111101","1000100011010011",
"0000110101000001","0001001000010001","0001000110000110","1000010010101111","1001010010011110","1001011010111000","1001001100100101","0001010001001100",
"0001100111011001","0001100111010010","0000110001001001","1001101101010111","1001110111100000","1001101101101111","0001100100000010","0010000001100100",
"0010000011001111","0001100011000110","1010000010110101","1010010001001000","1010001001010101","0001110001010100","0010010111100111","0010011101011001",
"0010000111000111","1010011000000000","1010101011000111","1010101001000001","0001110110101001","0010111001111100","0011001010001010","0011010001010110"
);

end FIR_Filter_2_package;

package body FIR_Filter_2_package is

end FIR_Filter_2_package;
